`default_nettype none
`timescale 1ns / 1ps

// module mem_cell #(parameter ADDR_BITS = 2) (
//   input clock,
//   input reset,
//   wire [ADDR_BITS-1:0] read_addr, write_addr,
//   wire we
// );
//   reg [7:0] mem[2**ADDR_BITS];

// endmodule